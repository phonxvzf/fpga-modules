`timescale 1ns / 1ns

module main(an, seg, dp, sw, clk);

output [3:0] an;
output [6:0] seg;
output reg dp = 0;
input wire [7:0] sw;
input wire clk;

endmodule
